--
--  Copyright 2011 Martin Schoeberl <masca@imm.dtu.dk>,
--                 Technical University of Denmark, DTU Informatics. 
--  All rights reserved.
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
-- 
--    1. Redistributions of source code must retain the above copyright notice,
--       this list of conditions and the following disclaimer.
-- 
--    2. Redistributions in binary form must reproduce the above copyright
--       notice, this list of conditions and the following disclaimer in the
--       documentation and/or other materials provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDER ``AS IS'' AND ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES
-- OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN
-- NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF
-- THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation are
-- those of the authors and should not be interpreted as representing official
-- policies, either expressed or implied, of the copyright holder.
-- 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

use work.leros_types.all;

-- instruction memory
-- write is ignored for now
-- the content should be generated by an assembler

entity leros_im is
	port  (
		clk : in std_logic;
		reset : in std_logic;
		din : in im_in_type;
		dout : out im_out_type
	);
end leros_im;

architecture rtl of leros_im is

	signal areg		: std_logic_vector(IM_BITS-1 downto 0);
	signal DOA		: std_logic_vector(31 downto 0);
	signal ADDRA   : std_logic_vector(13 downto 0);
	
	signal gndv    : std_logic_vector(31 downto 0);
	signal vccv    : std_logic_vector(15 downto 0);

begin

gndv <= "00000000000000000000000000000000";
vccv <= "1111111111111111";

process(clk) begin

	if rising_edge(clk) then
		areg <= din.rdaddr after 100 ps;
	end if;

end process;

	dout.data <= DOA(15 downto 0) after 100 ps;
	
	ADDRA <= din.rdaddr & "0000" after 100 ps;
	
	--rom: entity work.leros_rom port map(areg, data);
	  -- RAMB16BWER: 16k-bit Data and 2k-bit Parity Configurable Synchronous Dual Port Block RAM with Optional Output Registers
   --             Spartan-6
   -- Xilinx HDL Language Template, version 13.2

   RAMB16BWER_inst : RAMB16BWER
   generic map (
      -- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
      DATA_WIDTH_A => 18,
      DATA_WIDTH_B => 18,
      -- DOA_REG/DOB_REG: Optional output register (0 or 1)
      DOA_REG => 0,
      DOB_REG => 0,
      -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
      EN_RSTRAM_A => TRUE,
      EN_RSTRAM_B => TRUE,
      -- INITP_00 to INITP_07: Initial memory contents.
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- INIT_00 to INIT_3F: Initial memory contents.
      INIT_00 => X"40010000212530002172400100002125300021654001000021253000214c0000",
      INIT_01 => X"210a4001000021253000210d400100002125300021734001000021253000216f",
      INIT_02 => X"000000004001000020013801200049fd000023013c0048dd4001000021253000",
      INIT_03 => X"300d20083033300e200d3033200b30350c33000000004b0a200d3033200b3035",
      INIT_04 => X"20330c353033301e4809200b3033200d303520330c353033301e200e3033200c",
      INIT_05 => X"30350c33000000004b0c200e3033480248ba200c303520330c35303330204809",
      INIT_06 => X"200c3033200e303520330c35303330203033000000004a0248ec201e30330000",
      INIT_07 => X"00004a0248e6200b3033200d30350c33000000004b0421ff3022480321013022",
      INIT_08 => X"200c3033200e30350c33000000004b0421ff3024480321013024201e30332020",
      INIT_09 => X"303520330c35000000004c58202030330833303330263033201e303508353035",
      INIT_0A => X"20330c353033302820263033201e303520330c353033300f201e303300000000",
      INIT_0B => X"4c6220093033480248a420333800200a30333800200b30333800200c30333800",
      INIT_0C => X"200b30332022303508333033300b200f3033000000004c094908200c30332024",
      INIT_0D => X"303508333033300c200f3033000000004c0a4909200f30332028303508333033",
      INIT_0E => X"300f4808200f30332026303508333033300f201e0d01301e48c0201e30330833",
      INIT_0F => X"303330263033202030350835303520330c353033302820263033202030352033",
      INIT_10 => X"0c353033300f20203033000000004c0b20093033480248a920333800200a3033",
      INIT_11 => X"3800200b30333800200c30333800200c30332024303508333033300c200f3033",
      INIT_12 => X"000000004c094908200b30332022303508333033300b200f3033000000004c0a",
      INIT_13 => X"4909200f30332028303508333033300f4808200f30332026303508333033300f",
      INIT_14 => X"20200d01302048c0000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- INIT_A/INIT_B: Initial values on output port
      INIT_A => X"000000000",
      INIT_B => X"000000000",
      -- INIT_FILE: Optional file used to specify initial RAM contents
      INIT_FILE => "NONE",
      -- RSTTYPE: "SYNC" or "ASYNC" 
      RSTTYPE => "SYNC",
      -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
      RST_PRIORITY_A => "CE",
      RST_PRIORITY_B => "CE",
      -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
      SIM_COLLISION_CHECK => "ALL",
      -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
      SIM_DEVICE => "SPARTAN6",
      -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
      SRVAL_A => X"000000000",
      SRVAL_B => X"000000000",
      -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST" 
   )
   port map (
      -- Port A Data: 32-bit (each) output: Port A data
      DOA => DOA,       -- 32-bit output: A port data output
  --    DOPA => DOPA,     -- 4-bit output: A port parity output
      -- Port B Data: 32-bit (each) output: Port B data
  --    DOB => DOB,       -- 32-bit output: B port data output
  --    DOPB => DOPB,     -- 4-bit output: B port parity output
      -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
      ADDRA => ADDRA,   -- 14-bit input: A port address input
      CLKA => clk,     -- 1-bit input: A port clock input
      ENA => vccv(0),       -- 1-bit input: A port enable input
      REGCEA => vccv(0), -- 1-bit input: A port register clock enable input
      RSTA => gndv(0),     -- 1-bit input: A port register set/reset input
      WEA => gndv(3 downto 0),       -- 4-bit input: Port A byte-wide write enable input
      -- Port A Data: 32-bit (each) input: Port A data
      DIA => gndv(31 downto 0),       -- 32-bit input: A port data input
      DIPA => gndv(3 downto 0),     -- 4-bit input: A port parity input
      -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
      ADDRB => gndv(13 downto 0),   -- 14-bit input: B port address input
      CLKB => gndv(0),     -- 1-bit input: B port clock input
      ENB => gndv(0),       -- 1-bit input: B port enable input
      REGCEB => gndv(0), -- 1-bit input: B port register clock enable input
      RSTB => gndv(0),     -- 1-bit input: B port register set/reset input
      WEB => gndv(3 downto 0),       -- 4-bit input: Port B byte-wide write enable input
      -- Port B Data: 32-bit (each) input: Port B data
      DIB => gndv(31 downto 0),       -- 32-bit input: B port data input
      DIPB => gndv(3 downto 0)      -- 4-bit input: B port parity input
   );

--	rom : imem port map(
--		clka => clk,
 --    wea => gndv(0 downto 0),
  --   addra => din.rdaddr, 
   --  dina => gndv, 
  --   douta =>data);
	
-- use generated table
-- process(areg) begin
-- 
-- 	case areg is
-- 
-- 		when X"00" => data <= X"0000"; -- never executed
-- 		when X"01" => data <= X"0805"; -- load imm
-- 		when X"02" => data <= X"0e01"; -- sub 1 
-- 		when X"03" => data <= X"0e01"; -- sub 1 
-- 		when X"04" => data <= X"f000"; -- nop
-- 		when X"05" => data <= X"10fe"; -- brnz
-- 		when X"06" => data <= X"f000"; -- nop
-- 		when X"07" => data <= X"0801"; -- load 1
-- 		when X"08" => data <= X"2000"; -- outp
-- 		when X"09" => data <= X"0805"; -- load imm
-- 		when X"0a" => data <= X"0e01"; -- sub 1 
-- 		when X"0b" => data <= X"0e01"; -- sub 1 
-- 		when X"0c" => data <= X"f000"; -- nop
-- 		when X"0d" => data <= X"10fe"; -- brnz
-- 		when X"0e" => data <= X"f000"; -- nop
-- 		when X"0f" => data <= X"0800"; -- load 0
-- 		when X"10" => data <= X"2000"; -- outp
-- 		when X"11" => data <= X"0801"; -- load imm
-- 		when X"12" => data <= X"f000"; -- nop
-- 		when X"13" => data <= X"10ee"; -- brnz
-- 		when others => data <= X"f000"; 
-- 	end case;
-- end process;

end rtl;
